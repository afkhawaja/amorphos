/*

Uses the OCL AXI-Lite interface to convert 32-bit PCI-e

*/

import AMITypes::*;

module DMA_PCIS_CONTROLLER(

);

endmodule
